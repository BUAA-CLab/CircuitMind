module opposite_number(
    input wire [7:0] in,
    output [7:0] out
);

    assign out = -in;

endmodule
