module not_gate_ref(
    input wire in,
    output wire out
);

assign out = ~in;

endmodule
